module MEM_WR_Reg();



endmodule 